// niosII.v

// Generated using ACDS version 15.0 153

`timescale 1 ps / 1 ps
module niosII (
		input  wire [3:0]  btn_export,                       //       btn.export
		input  wire        clk_clk,                          //       clk.clk
		output wire [22:0] flash_bus_tcm_address_out,        // flash_bus.tcm_address_out
		output wire [0:0]  flash_bus_tcm_outputenable_n_out, //          .tcm_outputenable_n_out
		output wire [0:0]  flash_bus_tcm_reset_n_out,        //          .tcm_reset_n_out
		output wire [0:0]  flash_bus_tcm_write_n_out,        //          .tcm_write_n_out
		inout  wire [7:0]  flash_bus_tcm_data_out,           //          .tcm_data_out
		output wire [0:0]  flash_bus_tcm_chipselect_n_out,   //          .tcm_chipselect_n_out
		output wire        gen_export,                       //       gen.export
		output wire [31:0] hex_export,                       //       hex.export
		output wire [7:0]  led_export,                       //       led.export
		output wire [20:0] ram_bus_tcm_address_out,          //   ram_bus.tcm_address_out
		output wire [1:0]  ram_bus_tcm_byteenable_n_out,     //          .tcm_byteenable_n_out
		output wire [0:0]  ram_bus_tcm_outputenable_n_out,   //          .tcm_outputenable_n_out
		output wire [0:0]  ram_bus_tcm_write_n_out,          //          .tcm_write_n_out
		inout  wire [15:0] ram_bus_tcm_data_out,             //          .tcm_data_out
		output wire [0:0]  ram_bus_tcm_chipselect_n_out,     //          .tcm_chipselect_n_out
		input  wire        reset_reset_n                     //     reset.reset_n
	);

	wire         ext_ram_ctl_tcm_data_outen;                                            // ext_ram_ctl:tcm_data_outen -> ext_ram_bus:tcs_tcm_data_outen
	wire         ext_ram_ctl_tcm_outputenable_n_out;                                    // ext_ram_ctl:tcm_outputenable_n_out -> ext_ram_bus:tcs_tcm_outputenable_n_out
	wire         ext_ram_ctl_tcm_request;                                               // ext_ram_ctl:tcm_request -> ext_ram_bus:request
	wire   [1:0] ext_ram_ctl_tcm_byteenable_n_out;                                      // ext_ram_ctl:tcm_byteenable_n_out -> ext_ram_bus:tcs_tcm_byteenable_n_out
	wire         ext_ram_ctl_tcm_write_n_out;                                           // ext_ram_ctl:tcm_write_n_out -> ext_ram_bus:tcs_tcm_write_n_out
	wire         ext_ram_ctl_tcm_grant;                                                 // ext_ram_bus:grant -> ext_ram_ctl:tcm_grant
	wire         ext_ram_ctl_tcm_chipselect_n_out;                                      // ext_ram_ctl:tcm_chipselect_n_out -> ext_ram_bus:tcs_tcm_chipselect_n_out
	wire  [20:0] ext_ram_ctl_tcm_address_out;                                           // ext_ram_ctl:tcm_address_out -> ext_ram_bus:tcs_tcm_address_out
	wire  [15:0] ext_ram_ctl_tcm_data_out;                                              // ext_ram_ctl:tcm_data_out -> ext_ram_bus:tcs_tcm_data_out
	wire  [15:0] ext_ram_ctl_tcm_data_in;                                               // ext_ram_bus:tcs_tcm_data_in -> ext_ram_ctl:tcm_data_in
	wire         ext_flash_ctl_tcm_data_outen;                                          // ext_flash_ctl:tcm_data_outen -> ext_flash_bus:tcs_tcm_data_outen
	wire         ext_flash_ctl_tcm_outputenable_n_out;                                  // ext_flash_ctl:tcm_outputenable_n_out -> ext_flash_bus:tcs_tcm_outputenable_n_out
	wire         ext_flash_ctl_tcm_request;                                             // ext_flash_ctl:tcm_request -> ext_flash_bus:request
	wire         ext_flash_ctl_tcm_write_n_out;                                         // ext_flash_ctl:tcm_write_n_out -> ext_flash_bus:tcs_tcm_write_n_out
	wire         ext_flash_ctl_tcm_grant;                                               // ext_flash_bus:grant -> ext_flash_ctl:tcm_grant
	wire         ext_flash_ctl_tcm_reset_n_out;                                         // ext_flash_ctl:tcm_reset_n_out -> ext_flash_bus:tcs_tcm_reset_n_out
	wire         ext_flash_ctl_tcm_chipselect_n_out;                                    // ext_flash_ctl:tcm_chipselect_n_out -> ext_flash_bus:tcs_tcm_chipselect_n_out
	wire  [22:0] ext_flash_ctl_tcm_address_out;                                         // ext_flash_ctl:tcm_address_out -> ext_flash_bus:tcs_tcm_address_out
	wire   [7:0] ext_flash_ctl_tcm_data_out;                                            // ext_flash_ctl:tcm_data_out -> ext_flash_bus:tcs_tcm_data_out
	wire   [7:0] ext_flash_ctl_tcm_data_in;                                             // ext_flash_bus:tcs_tcm_data_in -> ext_flash_ctl:tcm_data_in
	wire  [31:0] cpu_custom_instruction_master_result;                                  // cpu_custom_instruction_master_translator:ci_slave_result -> cpu:E_ci_combo_result
	wire         cpu_custom_instruction_master_readra;                                  // cpu:E_ci_combo_readra -> cpu_custom_instruction_master_translator:ci_slave_readra
	wire   [4:0] cpu_custom_instruction_master_a;                                       // cpu:E_ci_combo_a -> cpu_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] cpu_custom_instruction_master_b;                                       // cpu:E_ci_combo_b -> cpu_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] cpu_custom_instruction_master_c;                                       // cpu:E_ci_combo_c -> cpu_custom_instruction_master_translator:ci_slave_c
	wire         cpu_custom_instruction_master_readrb;                                  // cpu:E_ci_combo_readrb -> cpu_custom_instruction_master_translator:ci_slave_readrb
	wire         cpu_custom_instruction_master_estatus;                                 // cpu:E_ci_combo_estatus -> cpu_custom_instruction_master_translator:ci_slave_estatus
	wire  [31:0] cpu_custom_instruction_master_ipending;                                // cpu:E_ci_combo_ipending -> cpu_custom_instruction_master_translator:ci_slave_ipending
	wire  [31:0] cpu_custom_instruction_master_datab;                                   // cpu:E_ci_combo_datab -> cpu_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] cpu_custom_instruction_master_dataa;                                   // cpu:E_ci_combo_dataa -> cpu_custom_instruction_master_translator:ci_slave_dataa
	wire         cpu_custom_instruction_master_writerc;                                 // cpu:E_ci_combo_writerc -> cpu_custom_instruction_master_translator:ci_slave_writerc
	wire   [7:0] cpu_custom_instruction_master_n;                                       // cpu:E_ci_combo_n -> cpu_custom_instruction_master_translator:ci_slave_n
	wire  [31:0] cpu_custom_instruction_master_translator_comb_ci_master_result;        // cpu_custom_instruction_master_comb_xconnect:ci_slave_result -> cpu_custom_instruction_master_translator:comb_ci_master_result
	wire         cpu_custom_instruction_master_translator_comb_ci_master_readra;        // cpu_custom_instruction_master_translator:comb_ci_master_readra -> cpu_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [4:0] cpu_custom_instruction_master_translator_comb_ci_master_a;             // cpu_custom_instruction_master_translator:comb_ci_master_a -> cpu_custom_instruction_master_comb_xconnect:ci_slave_a
	wire   [4:0] cpu_custom_instruction_master_translator_comb_ci_master_b;             // cpu_custom_instruction_master_translator:comb_ci_master_b -> cpu_custom_instruction_master_comb_xconnect:ci_slave_b
	wire         cpu_custom_instruction_master_translator_comb_ci_master_readrb;        // cpu_custom_instruction_master_translator:comb_ci_master_readrb -> cpu_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire   [4:0] cpu_custom_instruction_master_translator_comb_ci_master_c;             // cpu_custom_instruction_master_translator:comb_ci_master_c -> cpu_custom_instruction_master_comb_xconnect:ci_slave_c
	wire         cpu_custom_instruction_master_translator_comb_ci_master_estatus;       // cpu_custom_instruction_master_translator:comb_ci_master_estatus -> cpu_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] cpu_custom_instruction_master_translator_comb_ci_master_ipending;      // cpu_custom_instruction_master_translator:comb_ci_master_ipending -> cpu_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire  [31:0] cpu_custom_instruction_master_translator_comb_ci_master_datab;         // cpu_custom_instruction_master_translator:comb_ci_master_datab -> cpu_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] cpu_custom_instruction_master_translator_comb_ci_master_dataa;         // cpu_custom_instruction_master_translator:comb_ci_master_dataa -> cpu_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire         cpu_custom_instruction_master_translator_comb_ci_master_writerc;       // cpu_custom_instruction_master_translator:comb_ci_master_writerc -> cpu_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire   [7:0] cpu_custom_instruction_master_translator_comb_ci_master_n;             // cpu_custom_instruction_master_translator:comb_ci_master_n -> cpu_custom_instruction_master_comb_xconnect:ci_slave_n
	wire  [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_result;         // cpu_custom_instruction_master_comb_slave_translator0:ci_slave_result -> cpu_custom_instruction_master_comb_xconnect:ci_master0_result
	wire         cpu_custom_instruction_master_comb_xconnect_ci_master0_readra;         // cpu_custom_instruction_master_comb_xconnect:ci_master0_readra -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [4:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_a;              // cpu_custom_instruction_master_comb_xconnect:ci_master0_a -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire   [4:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_b;              // cpu_custom_instruction_master_comb_xconnect:ci_master0_b -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire         cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb;         // cpu_custom_instruction_master_comb_xconnect:ci_master0_readrb -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire   [4:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_c;              // cpu_custom_instruction_master_comb_xconnect:ci_master0_c -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire         cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus;        // cpu_custom_instruction_master_comb_xconnect:ci_master0_estatus -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending;       // cpu_custom_instruction_master_comb_xconnect:ci_master0_ipending -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire  [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_datab;          // cpu_custom_instruction_master_comb_xconnect:ci_master0_datab -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa;          // cpu_custom_instruction_master_comb_xconnect:ci_master0_dataa -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire         cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc;        // cpu_custom_instruction_master_comb_xconnect:ci_master0_writerc -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire   [7:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_n;              // cpu_custom_instruction_master_comb_xconnect:ci_master0_n -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire  [31:0] cpu_custom_instruction_master_comb_slave_translator0_ci_master_result; // countones:ones -> cpu_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa;  // cpu_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> countones:din
	wire  [31:0] cpu_data_master_readdata;                                              // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                           // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                           // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [25:0] cpu_data_master_address;                                               // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                            // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                                  // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                                         // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                                 // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                             // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                                       // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                                    // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [24:0] cpu_instruction_master_address;                                        // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                           // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                                  // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;             // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                 // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_sigmadelta_0_avalon_slave_0_chipselect;              // mm_interconnect_0:sigmadelta_0_avalon_slave_0_chipselect -> sigmadelta_0:cs
	wire         mm_interconnect_0_sigmadelta_0_avalon_slave_0_write;                   // mm_interconnect_0:sigmadelta_0_avalon_slave_0_write -> sigmadelta_0:wr_n
	wire  [31:0] mm_interconnect_0_sigmadelta_0_avalon_slave_0_writedata;               // mm_interconnect_0:sigmadelta_0_avalon_slave_0_writedata -> sigmadelta_0:wr_data
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                        // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                         // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_performance_counter_0_control_slave_readdata;        // performance_counter_0:readdata -> mm_interconnect_0:performance_counter_0_control_slave_readdata
	wire   [3:0] mm_interconnect_0_performance_counter_0_control_slave_address;         // mm_interconnect_0:performance_counter_0_control_slave_address -> performance_counter_0:address
	wire         mm_interconnect_0_performance_counter_0_control_slave_begintransfer;   // mm_interconnect_0:performance_counter_0_control_slave_begintransfer -> performance_counter_0:begintransfer
	wire         mm_interconnect_0_performance_counter_0_control_slave_write;           // mm_interconnect_0:performance_counter_0_control_slave_write -> performance_counter_0:write
	wire  [31:0] mm_interconnect_0_performance_counter_0_control_slave_writedata;       // mm_interconnect_0:performance_counter_0_control_slave_writedata -> performance_counter_0:writedata
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;                      // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;                   // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;                   // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;                       // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                          // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;                    // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;                         // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;                     // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire         mm_interconnect_0_seven_seg_s1_chipselect;                             // mm_interconnect_0:seven_seg_s1_chipselect -> seven_seg:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_s1_readdata;                               // seven_seg:readdata -> mm_interconnect_0:seven_seg_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_s1_address;                                // mm_interconnect_0:seven_seg_s1_address -> seven_seg:address
	wire         mm_interconnect_0_seven_seg_s1_write;                                  // mm_interconnect_0:seven_seg_s1_write -> seven_seg:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_s1_writedata;                              // mm_interconnect_0:seven_seg_s1_writedata -> seven_seg:writedata
	wire         mm_interconnect_0_buttons_s1_chipselect;                               // mm_interconnect_0:buttons_s1_chipselect -> buttons:chipselect
	wire  [31:0] mm_interconnect_0_buttons_s1_readdata;                                 // buttons:readdata -> mm_interconnect_0:buttons_s1_readdata
	wire   [1:0] mm_interconnect_0_buttons_s1_address;                                  // mm_interconnect_0:buttons_s1_address -> buttons:address
	wire         mm_interconnect_0_buttons_s1_write;                                    // mm_interconnect_0:buttons_s1_write -> buttons:write_n
	wire  [31:0] mm_interconnect_0_buttons_s1_writedata;                                // mm_interconnect_0:buttons_s1_writedata -> buttons:writedata
	wire         mm_interconnect_0_sys_clk_timer_s1_chipselect;                         // mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_readdata;                           // sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_clk_timer_s1_address;                            // mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_0_sys_clk_timer_s1_write;                              // mm_interconnect_0:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_writedata;                          // mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire         mm_interconnect_0_high_res_timer_s1_chipselect;                        // mm_interconnect_0:high_res_timer_s1_chipselect -> high_res_timer:chipselect
	wire  [15:0] mm_interconnect_0_high_res_timer_s1_readdata;                          // high_res_timer:readdata -> mm_interconnect_0:high_res_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_high_res_timer_s1_address;                           // mm_interconnect_0:high_res_timer_s1_address -> high_res_timer:address
	wire         mm_interconnect_0_high_res_timer_s1_write;                             // mm_interconnect_0:high_res_timer_s1_write -> high_res_timer:write_n
	wire  [15:0] mm_interconnect_0_high_res_timer_s1_writedata;                         // mm_interconnect_0:high_res_timer_s1_writedata -> high_res_timer:writedata
	wire         mm_interconnect_0_green_led_s1_chipselect;                             // mm_interconnect_0:green_led_s1_chipselect -> green_led:chipselect
	wire  [31:0] mm_interconnect_0_green_led_s1_readdata;                               // green_led:readdata -> mm_interconnect_0:green_led_s1_readdata
	wire   [1:0] mm_interconnect_0_green_led_s1_address;                                // mm_interconnect_0:green_led_s1_address -> green_led:address
	wire         mm_interconnect_0_green_led_s1_write;                                  // mm_interconnect_0:green_led_s1_write -> green_led:write_n
	wire  [31:0] mm_interconnect_0_green_led_s1_writedata;                              // mm_interconnect_0:green_led_s1_writedata -> green_led:writedata
	wire         mm_interconnect_0_instruction_tcm_s2_chipselect;                       // mm_interconnect_0:instruction_tcm_s2_chipselect -> instruction_tcm:chipselect2
	wire  [31:0] mm_interconnect_0_instruction_tcm_s2_readdata;                         // instruction_tcm:readdata2 -> mm_interconnect_0:instruction_tcm_s2_readdata
	wire  [11:0] mm_interconnect_0_instruction_tcm_s2_address;                          // mm_interconnect_0:instruction_tcm_s2_address -> instruction_tcm:address2
	wire   [3:0] mm_interconnect_0_instruction_tcm_s2_byteenable;                       // mm_interconnect_0:instruction_tcm_s2_byteenable -> instruction_tcm:byteenable2
	wire         mm_interconnect_0_instruction_tcm_s2_write;                            // mm_interconnect_0:instruction_tcm_s2_write -> instruction_tcm:write2
	wire  [31:0] mm_interconnect_0_instruction_tcm_s2_writedata;                        // mm_interconnect_0:instruction_tcm_s2_writedata -> instruction_tcm:writedata2
	wire         mm_interconnect_0_instruction_tcm_s2_clken;                            // mm_interconnect_0:instruction_tcm_s2_clken -> instruction_tcm:clken2
	wire  [15:0] mm_interconnect_0_ext_ram_ctl_uas_readdata;                            // ext_ram_ctl:uas_readdata -> mm_interconnect_0:ext_ram_ctl_uas_readdata
	wire         mm_interconnect_0_ext_ram_ctl_uas_waitrequest;                         // ext_ram_ctl:uas_waitrequest -> mm_interconnect_0:ext_ram_ctl_uas_waitrequest
	wire         mm_interconnect_0_ext_ram_ctl_uas_debugaccess;                         // mm_interconnect_0:ext_ram_ctl_uas_debugaccess -> ext_ram_ctl:uas_debugaccess
	wire  [20:0] mm_interconnect_0_ext_ram_ctl_uas_address;                             // mm_interconnect_0:ext_ram_ctl_uas_address -> ext_ram_ctl:uas_address
	wire         mm_interconnect_0_ext_ram_ctl_uas_read;                                // mm_interconnect_0:ext_ram_ctl_uas_read -> ext_ram_ctl:uas_read
	wire   [1:0] mm_interconnect_0_ext_ram_ctl_uas_byteenable;                          // mm_interconnect_0:ext_ram_ctl_uas_byteenable -> ext_ram_ctl:uas_byteenable
	wire         mm_interconnect_0_ext_ram_ctl_uas_readdatavalid;                       // ext_ram_ctl:uas_readdatavalid -> mm_interconnect_0:ext_ram_ctl_uas_readdatavalid
	wire         mm_interconnect_0_ext_ram_ctl_uas_lock;                                // mm_interconnect_0:ext_ram_ctl_uas_lock -> ext_ram_ctl:uas_lock
	wire         mm_interconnect_0_ext_ram_ctl_uas_write;                               // mm_interconnect_0:ext_ram_ctl_uas_write -> ext_ram_ctl:uas_write
	wire  [15:0] mm_interconnect_0_ext_ram_ctl_uas_writedata;                           // mm_interconnect_0:ext_ram_ctl_uas_writedata -> ext_ram_ctl:uas_writedata
	wire   [1:0] mm_interconnect_0_ext_ram_ctl_uas_burstcount;                          // mm_interconnect_0:ext_ram_ctl_uas_burstcount -> ext_ram_ctl:uas_burstcount
	wire   [7:0] mm_interconnect_0_ext_flash_ctl_uas_readdata;                          // ext_flash_ctl:uas_readdata -> mm_interconnect_0:ext_flash_ctl_uas_readdata
	wire         mm_interconnect_0_ext_flash_ctl_uas_waitrequest;                       // ext_flash_ctl:uas_waitrequest -> mm_interconnect_0:ext_flash_ctl_uas_waitrequest
	wire         mm_interconnect_0_ext_flash_ctl_uas_debugaccess;                       // mm_interconnect_0:ext_flash_ctl_uas_debugaccess -> ext_flash_ctl:uas_debugaccess
	wire  [22:0] mm_interconnect_0_ext_flash_ctl_uas_address;                           // mm_interconnect_0:ext_flash_ctl_uas_address -> ext_flash_ctl:uas_address
	wire         mm_interconnect_0_ext_flash_ctl_uas_read;                              // mm_interconnect_0:ext_flash_ctl_uas_read -> ext_flash_ctl:uas_read
	wire   [0:0] mm_interconnect_0_ext_flash_ctl_uas_byteenable;                        // mm_interconnect_0:ext_flash_ctl_uas_byteenable -> ext_flash_ctl:uas_byteenable
	wire         mm_interconnect_0_ext_flash_ctl_uas_readdatavalid;                     // ext_flash_ctl:uas_readdatavalid -> mm_interconnect_0:ext_flash_ctl_uas_readdatavalid
	wire         mm_interconnect_0_ext_flash_ctl_uas_lock;                              // mm_interconnect_0:ext_flash_ctl_uas_lock -> ext_flash_ctl:uas_lock
	wire         mm_interconnect_0_ext_flash_ctl_uas_write;                             // mm_interconnect_0:ext_flash_ctl_uas_write -> ext_flash_ctl:uas_write
	wire   [7:0] mm_interconnect_0_ext_flash_ctl_uas_writedata;                         // mm_interconnect_0:ext_flash_ctl_uas_writedata -> ext_flash_ctl:uas_writedata
	wire   [0:0] mm_interconnect_0_ext_flash_ctl_uas_burstcount;                        // mm_interconnect_0:ext_flash_ctl_uas_burstcount -> ext_flash_ctl:uas_burstcount
	wire  [31:0] cpu_tightly_coupled_instruction_master_0_readdata;                     // mm_interconnect_1:cpu_tightly_coupled_instruction_master_0_readdata -> cpu:icm0_readdata
	wire         cpu_tightly_coupled_instruction_master_0_waitrequest;                  // mm_interconnect_1:cpu_tightly_coupled_instruction_master_0_waitrequest -> cpu:icm0_waitrequest
	wire  [25:0] cpu_tightly_coupled_instruction_master_0_address;                      // cpu:icm0_address -> mm_interconnect_1:cpu_tightly_coupled_instruction_master_0_address
	wire         cpu_tightly_coupled_instruction_master_0_read;                         // cpu:icm0_read -> mm_interconnect_1:cpu_tightly_coupled_instruction_master_0_read
	wire         cpu_tightly_coupled_instruction_master_0_readdatavalid;                // mm_interconnect_1:cpu_tightly_coupled_instruction_master_0_readdatavalid -> cpu:icm0_readdatavalid
	wire         cpu_tightly_coupled_instruction_master_0_clken;                        // cpu:icm0_clken -> mm_interconnect_1:cpu_tightly_coupled_instruction_master_0_clken
	wire         mm_interconnect_1_instruction_tcm_s1_chipselect;                       // mm_interconnect_1:instruction_tcm_s1_chipselect -> instruction_tcm:chipselect
	wire  [31:0] mm_interconnect_1_instruction_tcm_s1_readdata;                         // instruction_tcm:readdata -> mm_interconnect_1:instruction_tcm_s1_readdata
	wire  [11:0] mm_interconnect_1_instruction_tcm_s1_address;                          // mm_interconnect_1:instruction_tcm_s1_address -> instruction_tcm:address
	wire   [3:0] mm_interconnect_1_instruction_tcm_s1_byteenable;                       // mm_interconnect_1:instruction_tcm_s1_byteenable -> instruction_tcm:byteenable
	wire         mm_interconnect_1_instruction_tcm_s1_write;                            // mm_interconnect_1:instruction_tcm_s1_write -> instruction_tcm:write
	wire  [31:0] mm_interconnect_1_instruction_tcm_s1_writedata;                        // mm_interconnect_1:instruction_tcm_s1_writedata -> instruction_tcm:writedata
	wire         mm_interconnect_1_instruction_tcm_s1_clken;                            // mm_interconnect_1:instruction_tcm_s1_clken -> instruction_tcm:clken
	wire         irq_mapper_receiver0_irq;                                              // sys_clk_timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                              // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                              // buttons:irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu_d_irq_irq;                                                         // irq_mapper:sender_irq -> cpu:d_irq
	wire         rst_controller_reset_out_reset;                                        // rst_controller:reset_out -> [buttons:reset_n, cpu:reset_n, ext_flash_bus:reset, ext_flash_ctl:reset_reset, ext_ram_bus:reset, ext_ram_ctl:reset_reset, green_led:reset_n, high_res_timer:reset_n, instruction_tcm:reset, instruction_tcm:reset2, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, mm_interconnect_1:cpu_reset_n_reset_bridge_in_reset_reset, performance_counter_0:reset_n, rst_translator:in_reset, seven_seg:reset_n, sigmadelta_0:clrn, sys_clk_timer:reset_n, sysid:reset_n]
	wire         rst_controller_reset_out_reset_req;                                    // rst_controller:reset_req -> [cpu:reset_req, instruction_tcm:reset_req, instruction_tcm:reset_req2, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                                     // cpu:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	niosII_buttons buttons (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_buttons_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_buttons_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_buttons_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_buttons_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_buttons_s1_readdata),   //                    .readdata
		.in_port    (btn_export),                              // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                 //                 irq.irq
	);

	countones countones (
		.din  (cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // nios_custom_instruction_slave.dataa
		.ones (cpu_custom_instruction_master_comb_slave_translator0_ci_master_result)  //                              .result
	);

	niosII_cpu cpu (
		.clk                                   (clk_clk),                                                //                                  clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                        //                              reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                     //                                     .reset_req
		.d_address                             (cpu_data_master_address),                                //                          data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                             //                                     .byteenable
		.d_read                                (cpu_data_master_read),                                   //                                     .read
		.d_readdata                            (cpu_data_master_readdata),                               //                                     .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                            //                                     .waitrequest
		.d_write                               (cpu_data_master_write),                                  //                                     .write
		.d_writedata                           (cpu_data_master_writedata),                              //                                     .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                          //                                     .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                            //                                     .debugaccess
		.i_address                             (cpu_instruction_master_address),                         //                   instruction_master.address
		.i_read                                (cpu_instruction_master_read),                            //                                     .read
		.i_readdata                            (cpu_instruction_master_readdata),                        //                                     .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                     //                                     .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                   //                                     .readdatavalid
		.icm0_readdata                         (cpu_tightly_coupled_instruction_master_0_readdata),      // tightly_coupled_instruction_master_0.readdata
		.icm0_waitrequest                      (cpu_tightly_coupled_instruction_master_0_waitrequest),   //                                     .waitrequest
		.icm0_readdatavalid                    (cpu_tightly_coupled_instruction_master_0_readdatavalid), //                                     .readdatavalid
		.icm0_address                          (cpu_tightly_coupled_instruction_master_0_address),       //                                     .address
		.icm0_read                             (cpu_tightly_coupled_instruction_master_0_read),          //                                     .read
		.icm0_clken                            (cpu_tightly_coupled_instruction_master_0_clken),         //                                     .clken
		.d_irq                                 (cpu_d_irq_irq),                                          //                                d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                      //              jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),        //                    jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),     //                                     .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),    //                                     .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),           //                                     .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),       //                                     .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),    //                                     .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),          //                                     .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),      //                                     .writedata
		.E_ci_combo_result                     (cpu_custom_instruction_master_result),                   //            custom_instruction_master.result
		.E_ci_combo_a                          (cpu_custom_instruction_master_a),                        //                                     .a
		.E_ci_combo_b                          (cpu_custom_instruction_master_b),                        //                                     .b
		.E_ci_combo_c                          (cpu_custom_instruction_master_c),                        //                                     .c
		.E_ci_combo_dataa                      (cpu_custom_instruction_master_dataa),                    //                                     .dataa
		.E_ci_combo_datab                      (cpu_custom_instruction_master_datab),                    //                                     .datab
		.E_ci_combo_estatus                    (cpu_custom_instruction_master_estatus),                  //                                     .estatus
		.E_ci_combo_ipending                   (cpu_custom_instruction_master_ipending),                 //                                     .ipending
		.E_ci_combo_n                          (cpu_custom_instruction_master_n),                        //                                     .n
		.E_ci_combo_readra                     (cpu_custom_instruction_master_readra),                   //                                     .readra
		.E_ci_combo_readrb                     (cpu_custom_instruction_master_readrb),                   //                                     .readrb
		.E_ci_combo_writerc                    (cpu_custom_instruction_master_writerc)                   //                                     .writerc
	);

	niosII_ext_flash_bus ext_flash_bus (
		.clk                        (clk_clk),                              //   clk.clk
		.reset                      (rst_controller_reset_out_reset),       // reset.reset
		.request                    (ext_flash_ctl_tcm_request),            //   tcs.request
		.grant                      (ext_flash_ctl_tcm_grant),              //      .grant
		.tcs_tcm_address_out        (ext_flash_ctl_tcm_address_out),        //      .address_out
		.tcs_tcm_outputenable_n_out (ext_flash_ctl_tcm_outputenable_n_out), //      .outputenable_n_out
		.tcs_tcm_reset_n_out        (ext_flash_ctl_tcm_reset_n_out),        //      .reset_n_out
		.tcs_tcm_write_n_out        (ext_flash_ctl_tcm_write_n_out),        //      .write_n_out
		.tcs_tcm_data_out           (ext_flash_ctl_tcm_data_out),           //      .data_out
		.tcs_tcm_data_outen         (ext_flash_ctl_tcm_data_outen),         //      .data_outen
		.tcs_tcm_data_in            (ext_flash_ctl_tcm_data_in),            //      .data_in
		.tcs_tcm_chipselect_n_out   (ext_flash_ctl_tcm_chipselect_n_out),   //      .chipselect_n_out
		.tcm_address_out            (flash_bus_tcm_address_out),            //   out.tcm_address_out
		.tcm_outputenable_n_out     (flash_bus_tcm_outputenable_n_out),     //      .tcm_outputenable_n_out
		.tcm_reset_n_out            (flash_bus_tcm_reset_n_out),            //      .tcm_reset_n_out
		.tcm_write_n_out            (flash_bus_tcm_write_n_out),            //      .tcm_write_n_out
		.tcm_data_out               (flash_bus_tcm_data_out),               //      .tcm_data_out
		.tcm_chipselect_n_out       (flash_bus_tcm_chipselect_n_out)        //      .tcm_chipselect_n_out
	);

	niosII_ext_flash_ctl #(
		.TCM_ADDRESS_W                  (23),
		.TCM_DATA_W                     (8),
		.TCM_BYTEENABLE_W               (1),
		.TCM_READ_WAIT                  (90),
		.TCM_WRITE_WAIT                 (90),
		.TCM_SETUP_WAIT                 (40),
		.TCM_DATA_HOLD                  (40),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (1),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (0),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (1),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (1),
		.ACTIVE_LOW_READ                (0),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (1),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) ext_flash_ctl (
		.clk_clk                (clk_clk),                                           //   clk.clk
		.reset_reset            (rst_controller_reset_out_reset),                    // reset.reset
		.uas_address            (mm_interconnect_0_ext_flash_ctl_uas_address),       //   uas.address
		.uas_burstcount         (mm_interconnect_0_ext_flash_ctl_uas_burstcount),    //      .burstcount
		.uas_read               (mm_interconnect_0_ext_flash_ctl_uas_read),          //      .read
		.uas_write              (mm_interconnect_0_ext_flash_ctl_uas_write),         //      .write
		.uas_waitrequest        (mm_interconnect_0_ext_flash_ctl_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid      (mm_interconnect_0_ext_flash_ctl_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable         (mm_interconnect_0_ext_flash_ctl_uas_byteenable),    //      .byteenable
		.uas_readdata           (mm_interconnect_0_ext_flash_ctl_uas_readdata),      //      .readdata
		.uas_writedata          (mm_interconnect_0_ext_flash_ctl_uas_writedata),     //      .writedata
		.uas_lock               (mm_interconnect_0_ext_flash_ctl_uas_lock),          //      .lock
		.uas_debugaccess        (mm_interconnect_0_ext_flash_ctl_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out        (ext_flash_ctl_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_chipselect_n_out   (ext_flash_ctl_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_outputenable_n_out (ext_flash_ctl_tcm_outputenable_n_out),              //      .outputenable_n_out
		.tcm_reset_n_out        (ext_flash_ctl_tcm_reset_n_out),                     //      .reset_n_out
		.tcm_request            (ext_flash_ctl_tcm_request),                         //      .request
		.tcm_grant              (ext_flash_ctl_tcm_grant),                           //      .grant
		.tcm_address_out        (ext_flash_ctl_tcm_address_out),                     //      .address_out
		.tcm_data_out           (ext_flash_ctl_tcm_data_out),                        //      .data_out
		.tcm_data_outen         (ext_flash_ctl_tcm_data_outen),                      //      .data_outen
		.tcm_data_in            (ext_flash_ctl_tcm_data_in)                          //      .data_in
	);

	niosII_ext_ram_bus ext_ram_bus (
		.clk                        (clk_clk),                            //   clk.clk
		.reset                      (rst_controller_reset_out_reset),     // reset.reset
		.request                    (ext_ram_ctl_tcm_request),            //   tcs.request
		.grant                      (ext_ram_ctl_tcm_grant),              //      .grant
		.tcs_tcm_address_out        (ext_ram_ctl_tcm_address_out),        //      .address_out
		.tcs_tcm_byteenable_n_out   (ext_ram_ctl_tcm_byteenable_n_out),   //      .byteenable_n_out
		.tcs_tcm_outputenable_n_out (ext_ram_ctl_tcm_outputenable_n_out), //      .outputenable_n_out
		.tcs_tcm_write_n_out        (ext_ram_ctl_tcm_write_n_out),        //      .write_n_out
		.tcs_tcm_data_out           (ext_ram_ctl_tcm_data_out),           //      .data_out
		.tcs_tcm_data_outen         (ext_ram_ctl_tcm_data_outen),         //      .data_outen
		.tcs_tcm_data_in            (ext_ram_ctl_tcm_data_in),            //      .data_in
		.tcs_tcm_chipselect_n_out   (ext_ram_ctl_tcm_chipselect_n_out),   //      .chipselect_n_out
		.tcm_address_out            (ram_bus_tcm_address_out),            //   out.tcm_address_out
		.tcm_byteenable_n_out       (ram_bus_tcm_byteenable_n_out),       //      .tcm_byteenable_n_out
		.tcm_outputenable_n_out     (ram_bus_tcm_outputenable_n_out),     //      .tcm_outputenable_n_out
		.tcm_write_n_out            (ram_bus_tcm_write_n_out),            //      .tcm_write_n_out
		.tcm_data_out               (ram_bus_tcm_data_out),               //      .tcm_data_out
		.tcm_chipselect_n_out       (ram_bus_tcm_chipselect_n_out)        //      .tcm_chipselect_n_out
	);

	niosII_ext_ram_ctl #(
		.TCM_ADDRESS_W                  (21),
		.TCM_DATA_W                     (16),
		.TCM_BYTEENABLE_W               (2),
		.TCM_READ_WAIT                  (20),
		.TCM_WRITE_WAIT                 (10),
		.TCM_SETUP_WAIT                 (5),
		.TCM_DATA_HOLD                  (10),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (2),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (0),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (1),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (1),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (0),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (1),
		.ACTIVE_LOW_OUTPUTENABLE        (1),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) ext_ram_ctl (
		.clk_clk                (clk_clk),                                         //   clk.clk
		.reset_reset            (rst_controller_reset_out_reset),                  // reset.reset
		.uas_address            (mm_interconnect_0_ext_ram_ctl_uas_address),       //   uas.address
		.uas_burstcount         (mm_interconnect_0_ext_ram_ctl_uas_burstcount),    //      .burstcount
		.uas_read               (mm_interconnect_0_ext_ram_ctl_uas_read),          //      .read
		.uas_write              (mm_interconnect_0_ext_ram_ctl_uas_write),         //      .write
		.uas_waitrequest        (mm_interconnect_0_ext_ram_ctl_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid      (mm_interconnect_0_ext_ram_ctl_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable         (mm_interconnect_0_ext_ram_ctl_uas_byteenable),    //      .byteenable
		.uas_readdata           (mm_interconnect_0_ext_ram_ctl_uas_readdata),      //      .readdata
		.uas_writedata          (mm_interconnect_0_ext_ram_ctl_uas_writedata),     //      .writedata
		.uas_lock               (mm_interconnect_0_ext_ram_ctl_uas_lock),          //      .lock
		.uas_debugaccess        (mm_interconnect_0_ext_ram_ctl_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out        (ext_ram_ctl_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_chipselect_n_out   (ext_ram_ctl_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_outputenable_n_out (ext_ram_ctl_tcm_outputenable_n_out),              //      .outputenable_n_out
		.tcm_request            (ext_ram_ctl_tcm_request),                         //      .request
		.tcm_grant              (ext_ram_ctl_tcm_grant),                           //      .grant
		.tcm_address_out        (ext_ram_ctl_tcm_address_out),                     //      .address_out
		.tcm_byteenable_n_out   (ext_ram_ctl_tcm_byteenable_n_out),                //      .byteenable_n_out
		.tcm_data_out           (ext_ram_ctl_tcm_data_out),                        //      .data_out
		.tcm_data_outen         (ext_ram_ctl_tcm_data_outen),                      //      .data_outen
		.tcm_data_in            (ext_ram_ctl_tcm_data_in)                          //      .data_in
	);

	niosII_green_led green_led (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_green_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_green_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_green_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_green_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_green_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                                 // external_connection.export
	);

	niosII_high_res_timer high_res_timer (
		.clk        (clk_clk),                                        //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                // reset.reset_n
		.address    (mm_interconnect_0_high_res_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_high_res_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_high_res_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_high_res_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_high_res_timer_s1_write),     //      .write_n
		.irq        ()                                                //   irq.irq
	);

	niosII_instruction_tcm instruction_tcm (
		.clk         (clk_clk),                                         //   clk1.clk
		.address     (mm_interconnect_1_instruction_tcm_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_instruction_tcm_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_instruction_tcm_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_instruction_tcm_s1_write),      //       .write
		.readdata    (mm_interconnect_1_instruction_tcm_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_instruction_tcm_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_1_instruction_tcm_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                  // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),              //       .reset_req
		.address2    (mm_interconnect_0_instruction_tcm_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_instruction_tcm_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_instruction_tcm_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_instruction_tcm_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_instruction_tcm_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_instruction_tcm_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_instruction_tcm_s2_byteenable), //       .byteenable
		.clk2        (clk_clk),                                         //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),                  // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req)               //       .reset_req
	);

	niosII_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	niosII_performance_counter_0 performance_counter_0 (
		.clk           (clk_clk),                                                             //           clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                     //         reset.reset_n
		.address       (mm_interconnect_0_performance_counter_0_control_slave_address),       // control_slave.address
		.begintransfer (mm_interconnect_0_performance_counter_0_control_slave_begintransfer), //              .begintransfer
		.readdata      (mm_interconnect_0_performance_counter_0_control_slave_readdata),      //              .readdata
		.write         (mm_interconnect_0_performance_counter_0_control_slave_write),         //              .write
		.writedata     (mm_interconnect_0_performance_counter_0_control_slave_writedata)      //              .writedata
	);

	niosII_seven_seg seven_seg (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_s1_readdata),   //                    .readdata
		.out_port   (hex_export)                                 // external_connection.export
	);

	sigmadelta sigmadelta_0 (
		.clk     (clk_clk),                                                  //          clock.clk
		.cs      (mm_interconnect_0_sigmadelta_0_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.wr_data (mm_interconnect_0_sigmadelta_0_avalon_slave_0_writedata),  //               .writedata
		.wr_n    (~mm_interconnect_0_sigmadelta_0_avalon_slave_0_write),     //               .write_n
		.clrn    (~rst_controller_reset_out_reset),                          //     reset_sink.reset_n
		.daco    (gen_export)                                                //    conduit_end.export
	);

	niosII_sys_clk_timer sys_clk_timer (
		.clk        (clk_clk),                                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                       //   irq.irq
	);

	niosII_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) cpu_custom_instruction_master_translator (
		.ci_slave_dataa            (cpu_custom_instruction_master_dataa),                              //       ci_slave.dataa
		.ci_slave_datab            (cpu_custom_instruction_master_datab),                              //               .datab
		.ci_slave_result           (cpu_custom_instruction_master_result),                             //               .result
		.ci_slave_n                (cpu_custom_instruction_master_n),                                  //               .n
		.ci_slave_readra           (cpu_custom_instruction_master_readra),                             //               .readra
		.ci_slave_readrb           (cpu_custom_instruction_master_readrb),                             //               .readrb
		.ci_slave_writerc          (cpu_custom_instruction_master_writerc),                            //               .writerc
		.ci_slave_a                (cpu_custom_instruction_master_a),                                  //               .a
		.ci_slave_b                (cpu_custom_instruction_master_b),                                  //               .b
		.ci_slave_c                (cpu_custom_instruction_master_c),                                  //               .c
		.ci_slave_ipending         (cpu_custom_instruction_master_ipending),                           //               .ipending
		.ci_slave_estatus          (cpu_custom_instruction_master_estatus),                            //               .estatus
		.comb_ci_master_dataa      (cpu_custom_instruction_master_translator_comb_ci_master_dataa),    // comb_ci_master.dataa
		.comb_ci_master_datab      (cpu_custom_instruction_master_translator_comb_ci_master_datab),    //               .datab
		.comb_ci_master_result     (cpu_custom_instruction_master_translator_comb_ci_master_result),   //               .result
		.comb_ci_master_n          (cpu_custom_instruction_master_translator_comb_ci_master_n),        //               .n
		.comb_ci_master_readra     (cpu_custom_instruction_master_translator_comb_ci_master_readra),   //               .readra
		.comb_ci_master_readrb     (cpu_custom_instruction_master_translator_comb_ci_master_readrb),   //               .readrb
		.comb_ci_master_writerc    (cpu_custom_instruction_master_translator_comb_ci_master_writerc),  //               .writerc
		.comb_ci_master_a          (cpu_custom_instruction_master_translator_comb_ci_master_a),        //               .a
		.comb_ci_master_b          (cpu_custom_instruction_master_translator_comb_ci_master_b),        //               .b
		.comb_ci_master_c          (cpu_custom_instruction_master_translator_comb_ci_master_c),        //               .c
		.comb_ci_master_ipending   (cpu_custom_instruction_master_translator_comb_ci_master_ipending), //               .ipending
		.comb_ci_master_estatus    (cpu_custom_instruction_master_translator_comb_ci_master_estatus),  //               .estatus
		.ci_slave_multi_clk        (1'b0),                                                             //    (terminated)
		.ci_slave_multi_reset      (1'b0),                                                             //    (terminated)
		.ci_slave_multi_clken      (1'b0),                                                             //    (terminated)
		.ci_slave_multi_reset_req  (1'b0),                                                             //    (terminated)
		.ci_slave_multi_start      (1'b0),                                                             //    (terminated)
		.ci_slave_multi_done       (),                                                                 //    (terminated)
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                             //    (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                             //    (terminated)
		.ci_slave_multi_result     (),                                                                 //    (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                      //    (terminated)
		.ci_slave_multi_readra     (1'b0),                                                             //    (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                             //    (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                             //    (terminated)
		.ci_slave_multi_a          (5'b00000),                                                         //    (terminated)
		.ci_slave_multi_b          (5'b00000),                                                         //    (terminated)
		.ci_slave_multi_c          (5'b00000),                                                         //    (terminated)
		.multi_ci_master_clk       (),                                                                 //    (terminated)
		.multi_ci_master_reset     (),                                                                 //    (terminated)
		.multi_ci_master_clken     (),                                                                 //    (terminated)
		.multi_ci_master_reset_req (),                                                                 //    (terminated)
		.multi_ci_master_start     (),                                                                 //    (terminated)
		.multi_ci_master_done      (1'b0),                                                             //    (terminated)
		.multi_ci_master_dataa     (),                                                                 //    (terminated)
		.multi_ci_master_datab     (),                                                                 //    (terminated)
		.multi_ci_master_result    (32'b00000000000000000000000000000000),                             //    (terminated)
		.multi_ci_master_n         (),                                                                 //    (terminated)
		.multi_ci_master_readra    (),                                                                 //    (terminated)
		.multi_ci_master_readrb    (),                                                                 //    (terminated)
		.multi_ci_master_writerc   (),                                                                 //    (terminated)
		.multi_ci_master_a         (),                                                                 //    (terminated)
		.multi_ci_master_b         (),                                                                 //    (terminated)
		.multi_ci_master_c         ()                                                                  //    (terminated)
	);

	niosII_cpu_custom_instruction_master_comb_xconnect cpu_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (cpu_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (cpu_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (cpu_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (cpu_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (cpu_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (cpu_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (cpu_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (cpu_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (cpu_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (cpu_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (cpu_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (cpu_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (cpu_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (cpu_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (cpu_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (cpu_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (cpu_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (cpu_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (cpu_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) cpu_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (cpu_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (cpu_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (cpu_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (cpu_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (cpu_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (cpu_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (cpu_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_result    (cpu_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_datab     (),                                                                      // (terminated)
		.ci_master_n         (),                                                                      // (terminated)
		.ci_master_readra    (),                                                                      // (terminated)
		.ci_master_readrb    (),                                                                      // (terminated)
		.ci_master_writerc   (),                                                                      // (terminated)
		.ci_master_a         (),                                                                      // (terminated)
		.ci_master_b         (),                                                                      // (terminated)
		.ci_master_c         (),                                                                      // (terminated)
		.ci_master_ipending  (),                                                                      // (terminated)
		.ci_master_estatus   (),                                                                      // (terminated)
		.ci_master_clk       (),                                                                      // (terminated)
		.ci_master_clken     (),                                                                      // (terminated)
		.ci_master_reset_req (),                                                                      // (terminated)
		.ci_master_reset     (),                                                                      // (terminated)
		.ci_master_start     (),                                                                      // (terminated)
		.ci_master_done      (1'b0),                                                                  // (terminated)
		.ci_slave_clk        (1'b0),                                                                  // (terminated)
		.ci_slave_clken      (1'b0),                                                                  // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                  // (terminated)
		.ci_slave_reset      (1'b0),                                                                  // (terminated)
		.ci_slave_start      (1'b0),                                                                  // (terminated)
		.ci_slave_done       ()                                                                       // (terminated)
	);

	niosII_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                       (clk_clk),                                                             //                             clk_clk.clk
		.cpu_reset_n_reset_bridge_in_reset_reset           (rst_controller_reset_out_reset),                                      //   cpu_reset_n_reset_bridge_in_reset.reset
		.cpu_data_master_address                           (cpu_data_master_address),                                             //                     cpu_data_master.address
		.cpu_data_master_waitrequest                       (cpu_data_master_waitrequest),                                         //                                    .waitrequest
		.cpu_data_master_byteenable                        (cpu_data_master_byteenable),                                          //                                    .byteenable
		.cpu_data_master_read                              (cpu_data_master_read),                                                //                                    .read
		.cpu_data_master_readdata                          (cpu_data_master_readdata),                                            //                                    .readdata
		.cpu_data_master_readdatavalid                     (cpu_data_master_readdatavalid),                                       //                                    .readdatavalid
		.cpu_data_master_write                             (cpu_data_master_write),                                               //                                    .write
		.cpu_data_master_writedata                         (cpu_data_master_writedata),                                           //                                    .writedata
		.cpu_data_master_debugaccess                       (cpu_data_master_debugaccess),                                         //                                    .debugaccess
		.cpu_instruction_master_address                    (cpu_instruction_master_address),                                      //              cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                (cpu_instruction_master_waitrequest),                                  //                                    .waitrequest
		.cpu_instruction_master_read                       (cpu_instruction_master_read),                                         //                                    .read
		.cpu_instruction_master_readdata                   (cpu_instruction_master_readdata),                                     //                                    .readdata
		.cpu_instruction_master_readdatavalid              (cpu_instruction_master_readdatavalid),                                //                                    .readdatavalid
		.buttons_s1_address                                (mm_interconnect_0_buttons_s1_address),                                //                          buttons_s1.address
		.buttons_s1_write                                  (mm_interconnect_0_buttons_s1_write),                                  //                                    .write
		.buttons_s1_readdata                               (mm_interconnect_0_buttons_s1_readdata),                               //                                    .readdata
		.buttons_s1_writedata                              (mm_interconnect_0_buttons_s1_writedata),                              //                                    .writedata
		.buttons_s1_chipselect                             (mm_interconnect_0_buttons_s1_chipselect),                             //                                    .chipselect
		.cpu_jtag_debug_module_address                     (mm_interconnect_0_cpu_jtag_debug_module_address),                     //               cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write                       (mm_interconnect_0_cpu_jtag_debug_module_write),                       //                                    .write
		.cpu_jtag_debug_module_read                        (mm_interconnect_0_cpu_jtag_debug_module_read),                        //                                    .read
		.cpu_jtag_debug_module_readdata                    (mm_interconnect_0_cpu_jtag_debug_module_readdata),                    //                                    .readdata
		.cpu_jtag_debug_module_writedata                   (mm_interconnect_0_cpu_jtag_debug_module_writedata),                   //                                    .writedata
		.cpu_jtag_debug_module_byteenable                  (mm_interconnect_0_cpu_jtag_debug_module_byteenable),                  //                                    .byteenable
		.cpu_jtag_debug_module_waitrequest                 (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),                 //                                    .waitrequest
		.cpu_jtag_debug_module_debugaccess                 (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),                 //                                    .debugaccess
		.ext_flash_ctl_uas_address                         (mm_interconnect_0_ext_flash_ctl_uas_address),                         //                   ext_flash_ctl_uas.address
		.ext_flash_ctl_uas_write                           (mm_interconnect_0_ext_flash_ctl_uas_write),                           //                                    .write
		.ext_flash_ctl_uas_read                            (mm_interconnect_0_ext_flash_ctl_uas_read),                            //                                    .read
		.ext_flash_ctl_uas_readdata                        (mm_interconnect_0_ext_flash_ctl_uas_readdata),                        //                                    .readdata
		.ext_flash_ctl_uas_writedata                       (mm_interconnect_0_ext_flash_ctl_uas_writedata),                       //                                    .writedata
		.ext_flash_ctl_uas_burstcount                      (mm_interconnect_0_ext_flash_ctl_uas_burstcount),                      //                                    .burstcount
		.ext_flash_ctl_uas_byteenable                      (mm_interconnect_0_ext_flash_ctl_uas_byteenable),                      //                                    .byteenable
		.ext_flash_ctl_uas_readdatavalid                   (mm_interconnect_0_ext_flash_ctl_uas_readdatavalid),                   //                                    .readdatavalid
		.ext_flash_ctl_uas_waitrequest                     (mm_interconnect_0_ext_flash_ctl_uas_waitrequest),                     //                                    .waitrequest
		.ext_flash_ctl_uas_lock                            (mm_interconnect_0_ext_flash_ctl_uas_lock),                            //                                    .lock
		.ext_flash_ctl_uas_debugaccess                     (mm_interconnect_0_ext_flash_ctl_uas_debugaccess),                     //                                    .debugaccess
		.ext_ram_ctl_uas_address                           (mm_interconnect_0_ext_ram_ctl_uas_address),                           //                     ext_ram_ctl_uas.address
		.ext_ram_ctl_uas_write                             (mm_interconnect_0_ext_ram_ctl_uas_write),                             //                                    .write
		.ext_ram_ctl_uas_read                              (mm_interconnect_0_ext_ram_ctl_uas_read),                              //                                    .read
		.ext_ram_ctl_uas_readdata                          (mm_interconnect_0_ext_ram_ctl_uas_readdata),                          //                                    .readdata
		.ext_ram_ctl_uas_writedata                         (mm_interconnect_0_ext_ram_ctl_uas_writedata),                         //                                    .writedata
		.ext_ram_ctl_uas_burstcount                        (mm_interconnect_0_ext_ram_ctl_uas_burstcount),                        //                                    .burstcount
		.ext_ram_ctl_uas_byteenable                        (mm_interconnect_0_ext_ram_ctl_uas_byteenable),                        //                                    .byteenable
		.ext_ram_ctl_uas_readdatavalid                     (mm_interconnect_0_ext_ram_ctl_uas_readdatavalid),                     //                                    .readdatavalid
		.ext_ram_ctl_uas_waitrequest                       (mm_interconnect_0_ext_ram_ctl_uas_waitrequest),                       //                                    .waitrequest
		.ext_ram_ctl_uas_lock                              (mm_interconnect_0_ext_ram_ctl_uas_lock),                              //                                    .lock
		.ext_ram_ctl_uas_debugaccess                       (mm_interconnect_0_ext_ram_ctl_uas_debugaccess),                       //                                    .debugaccess
		.green_led_s1_address                              (mm_interconnect_0_green_led_s1_address),                              //                        green_led_s1.address
		.green_led_s1_write                                (mm_interconnect_0_green_led_s1_write),                                //                                    .write
		.green_led_s1_readdata                             (mm_interconnect_0_green_led_s1_readdata),                             //                                    .readdata
		.green_led_s1_writedata                            (mm_interconnect_0_green_led_s1_writedata),                            //                                    .writedata
		.green_led_s1_chipselect                           (mm_interconnect_0_green_led_s1_chipselect),                           //                                    .chipselect
		.high_res_timer_s1_address                         (mm_interconnect_0_high_res_timer_s1_address),                         //                   high_res_timer_s1.address
		.high_res_timer_s1_write                           (mm_interconnect_0_high_res_timer_s1_write),                           //                                    .write
		.high_res_timer_s1_readdata                        (mm_interconnect_0_high_res_timer_s1_readdata),                        //                                    .readdata
		.high_res_timer_s1_writedata                       (mm_interconnect_0_high_res_timer_s1_writedata),                       //                                    .writedata
		.high_res_timer_s1_chipselect                      (mm_interconnect_0_high_res_timer_s1_chipselect),                      //                                    .chipselect
		.instruction_tcm_s2_address                        (mm_interconnect_0_instruction_tcm_s2_address),                        //                  instruction_tcm_s2.address
		.instruction_tcm_s2_write                          (mm_interconnect_0_instruction_tcm_s2_write),                          //                                    .write
		.instruction_tcm_s2_readdata                       (mm_interconnect_0_instruction_tcm_s2_readdata),                       //                                    .readdata
		.instruction_tcm_s2_writedata                      (mm_interconnect_0_instruction_tcm_s2_writedata),                      //                                    .writedata
		.instruction_tcm_s2_byteenable                     (mm_interconnect_0_instruction_tcm_s2_byteenable),                     //                                    .byteenable
		.instruction_tcm_s2_chipselect                     (mm_interconnect_0_instruction_tcm_s2_chipselect),                     //                                    .chipselect
		.instruction_tcm_s2_clken                          (mm_interconnect_0_instruction_tcm_s2_clken),                          //                                    .clken
		.jtag_uart_avalon_jtag_slave_address               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),               //         jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                 //                                    .write
		.jtag_uart_avalon_jtag_slave_read                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                  //                                    .read
		.jtag_uart_avalon_jtag_slave_readdata              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),              //                                    .readdata
		.jtag_uart_avalon_jtag_slave_writedata             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),             //                                    .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),           //                                    .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),            //                                    .chipselect
		.performance_counter_0_control_slave_address       (mm_interconnect_0_performance_counter_0_control_slave_address),       // performance_counter_0_control_slave.address
		.performance_counter_0_control_slave_write         (mm_interconnect_0_performance_counter_0_control_slave_write),         //                                    .write
		.performance_counter_0_control_slave_readdata      (mm_interconnect_0_performance_counter_0_control_slave_readdata),      //                                    .readdata
		.performance_counter_0_control_slave_writedata     (mm_interconnect_0_performance_counter_0_control_slave_writedata),     //                                    .writedata
		.performance_counter_0_control_slave_begintransfer (mm_interconnect_0_performance_counter_0_control_slave_begintransfer), //                                    .begintransfer
		.seven_seg_s1_address                              (mm_interconnect_0_seven_seg_s1_address),                              //                        seven_seg_s1.address
		.seven_seg_s1_write                                (mm_interconnect_0_seven_seg_s1_write),                                //                                    .write
		.seven_seg_s1_readdata                             (mm_interconnect_0_seven_seg_s1_readdata),                             //                                    .readdata
		.seven_seg_s1_writedata                            (mm_interconnect_0_seven_seg_s1_writedata),                            //                                    .writedata
		.seven_seg_s1_chipselect                           (mm_interconnect_0_seven_seg_s1_chipselect),                           //                                    .chipselect
		.sigmadelta_0_avalon_slave_0_write                 (mm_interconnect_0_sigmadelta_0_avalon_slave_0_write),                 //         sigmadelta_0_avalon_slave_0.write
		.sigmadelta_0_avalon_slave_0_writedata             (mm_interconnect_0_sigmadelta_0_avalon_slave_0_writedata),             //                                    .writedata
		.sigmadelta_0_avalon_slave_0_chipselect            (mm_interconnect_0_sigmadelta_0_avalon_slave_0_chipselect),            //                                    .chipselect
		.sys_clk_timer_s1_address                          (mm_interconnect_0_sys_clk_timer_s1_address),                          //                    sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                            (mm_interconnect_0_sys_clk_timer_s1_write),                            //                                    .write
		.sys_clk_timer_s1_readdata                         (mm_interconnect_0_sys_clk_timer_s1_readdata),                         //                                    .readdata
		.sys_clk_timer_s1_writedata                        (mm_interconnect_0_sys_clk_timer_s1_writedata),                        //                                    .writedata
		.sys_clk_timer_s1_chipselect                       (mm_interconnect_0_sys_clk_timer_s1_chipselect),                       //                                    .chipselect
		.sysid_control_slave_address                       (mm_interconnect_0_sysid_control_slave_address),                       //                 sysid_control_slave.address
		.sysid_control_slave_readdata                      (mm_interconnect_0_sysid_control_slave_readdata)                       //                                    .readdata
	);

	niosII_mm_interconnect_1 mm_interconnect_1 (
		.clk_clk_clk                                            (clk_clk),                                                //                                  clk_clk.clk
		.cpu_reset_n_reset_bridge_in_reset_reset                (rst_controller_reset_out_reset),                         //        cpu_reset_n_reset_bridge_in_reset.reset
		.cpu_tightly_coupled_instruction_master_0_address       (cpu_tightly_coupled_instruction_master_0_address),       // cpu_tightly_coupled_instruction_master_0.address
		.cpu_tightly_coupled_instruction_master_0_waitrequest   (cpu_tightly_coupled_instruction_master_0_waitrequest),   //                                         .waitrequest
		.cpu_tightly_coupled_instruction_master_0_read          (cpu_tightly_coupled_instruction_master_0_read),          //                                         .read
		.cpu_tightly_coupled_instruction_master_0_readdata      (cpu_tightly_coupled_instruction_master_0_readdata),      //                                         .readdata
		.cpu_tightly_coupled_instruction_master_0_readdatavalid (cpu_tightly_coupled_instruction_master_0_readdatavalid), //                                         .readdatavalid
		.cpu_tightly_coupled_instruction_master_0_clken         (cpu_tightly_coupled_instruction_master_0_clken),         //                                         .clken
		.instruction_tcm_s1_address                             (mm_interconnect_1_instruction_tcm_s1_address),           //                       instruction_tcm_s1.address
		.instruction_tcm_s1_write                               (mm_interconnect_1_instruction_tcm_s1_write),             //                                         .write
		.instruction_tcm_s1_readdata                            (mm_interconnect_1_instruction_tcm_s1_readdata),          //                                         .readdata
		.instruction_tcm_s1_writedata                           (mm_interconnect_1_instruction_tcm_s1_writedata),         //                                         .writedata
		.instruction_tcm_s1_byteenable                          (mm_interconnect_1_instruction_tcm_s1_byteenable),        //                                         .byteenable
		.instruction_tcm_s1_chipselect                          (mm_interconnect_1_instruction_tcm_s1_chipselect),        //                                         .chipselect
		.instruction_tcm_s1_clken                               (mm_interconnect_1_instruction_tcm_s1_clken)              //                                         .clken
	);

	niosII_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
